package definitions;
parameter int CLOCK_PERIOD = 100; // 10 MHz
endpackage