//////////////////////////////////////////////////////////////////////////////////                                                           
// Third Year Project: RISC-V RV32i Pipelined Processor
// File: Writeback                                                   
// Description: Holds all Writeback stage modules.
//              Data Memory: 
//                  Holds the data for the program to operate on and allows read/writes. Follows a single-port BRAM template.
// Author: Luke Shepherd
// Date Modified: February 2025                                                                                                                                                                                                                                                       
//////////////////////////////////////////////////////////////////////////////////

module writeback ();
endmodule