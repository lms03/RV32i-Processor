//////////////////////////////////////////////////////////////////////////////////                                                           
// Third Year Project: RISC-V RV32i Pipelined Processor
// File: Extender                                                   
// Description: Generic extender used to sign extend the immediate and sign/zero extend loaded bytes/halfwords.
// Author: Luke Shepherd                                                     
// Date Created: November 2024                                                                                                                                                                                                                                                       
//////////////////////////////////////////////////////////////////////////////////

module extender (

);
endmodule